library verilog;
use verilog.vl_types.all;
entity mips_data_mem_testbench is
end mips_data_mem_testbench;
