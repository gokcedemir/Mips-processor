library verilog;
use verilog.vl_types.all;
entity mips_inst_mem_testbench is
end mips_inst_mem_testbench;
